// 2x2ConvTree GENERATED FROM CADA but shifter to upper right of compute array so fits in with 3x3ConvTree.
// This TB to get correct latency aligned for 2x2 convolutions kernels for layer 2.

`timescale 1ns / 1ns

module K3_E216B_2x2ConvTree_upperRight_layer2_latencyTest_RTL_TB();
reg  clk, rst; 
wire [143:0] dataOut; 
reg [1727:0] dataIn; 
reg [6:0] configIn; 
reg [35:0] controlIn; 
reg [125:0] gcontrolIn; 
reg [15:0] selectedChannel; 

// To test latency of inputs of layer2 with 2x2 kernel of stride 2.
reg [255:0] L2in; // Layer 2 input = input to 2x2 convolution with stride = 2.
reg [63:0] K2;  //  Layer 2 2x2 convolution kernel

ArrayTop uut(
.clk(clk),
.rst(rst),
.dataOut(dataOut),
.dataIn(dataIn),
.configIn(configIn),
.controlIn(controlIn),
.gControlIn(gcontrolIn)
);

always #1 clk = ~clk;

initial begin;

rst = 1'b1;
clk = 1'b1;
dataIn = 0;

L2in = {
16'd156,  16'd192,  16'd228,  16'd264,
16'd192,  16'd228,  16'd264,  16'd300,
16'd228,  16'd264,  16'd300,  16'd336,
16'd264,  16'd300,  16'd336,  16'd372 };

K2 = {
16'd2,  16'd3,
16'd3,  16'd4 };

#20
rst = 1'b0;
// Send in configuration bitstream - SHIFTED ALL controlIn bits to the right by 4 so 2x2convTree fits in upper right corner of array.
configIn =7'b0000000; 
controlIn =36'b000010000000000000000000000000000000;    // 1's shifted 4 bits over.
#2
configIn =7'b1101000; 
controlIn =36'b000001000000000000000000000000000000;    // 1's shifted 4 bits over. 
#2
configIn =7'b0000001; 
controlIn =36'b000000000000000011000000000000000000;    // 1's shifted 4 bits over. 
#2
configIn =7'b0100010; 
controlIn =36'b000000000011000000000000000000000000;    // 1's shifted 4 bits over. 
#2

// !!ORIGINAL!! This is your output channel 
// assign selectedChannel =  dataOut[15:0]; 
// !!NEW!! Shifted over by 2 output channels. This is your output channel 
assign selectedChannel =  dataOut[47:32];

// !!ORIGINAL!! Your input IO Config
//000000000000000000000000000000000000000000000000000000000000000000110110000000000000110110000000000000000000
// !!NEW!! Shifted 12 bits to the left. Your input IO Config
//000000000000000000000000000000000000000000000000000000110110000000000000110110000000000000000000000000000000

// !!ORIGINAL!! Your output IO Config
//000000000000000001
// !!ORIGINAL!! Your output IO Config
//000000000000010000
// Put together
// !!ORIGINAL!! Send in IO Configuration 
//gcontrolIn =126'b000000000000000001000000000000000000000000000000000000000000000000000000000000000000110110000000000000110110000000000000000000; 
// !!NEW!! Send in IO Configuration 
gcontrolIn =126'b000000000000010000000000000000000000000000000000000000000000000000000000110110000000000000110110000000000000000000000000000000; 
#2

/* // !!ORIGINAL!! 2x2convTree INPUT MAP ('IN1' to 'IN8'). Maps to 'Your input IO Config' 1 locations above.
dataIn = {
16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  IN7,IN8,16'd0,      IN3,IN4,16'd0,  
16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  IN5,IN6,16'd0,      IN1,IN2,16'd0,  
16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0};
*/

/* // !!NEW!! 2x2convTree INPUT MAP + LATENCY ('IN1_Lx' to 'IN8_Lx'). Maps to 'Your input IO Config' 1 locations above.
dataIn = {
16'd0,16'd0,16'd0,      16'd0,16'd0,16'd0,      16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
16'd0,16'd0,16'd0,      16'd0,16'd0,16'd0,      16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
16'd0,16'd0,16'd0,      16'd0,16'd0,16'd0,      16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
IN7_L1,IN8_L1,16'd0,    IN3_L2,IN4_L1,16'd0,    16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
IN5_L2,IN6_L2,16'd0,    IN1_L2,IN2_L2,16'd0,    16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
16'd0,16'd0,16'd0,      16'd0,16'd0,16'd0,      16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0};

  "inputLatency": [
      2,
      2,
      1,
      1,
      2,
      2,
      1,
      1
  ],
  
  Inputs 1, 2, 5 and 6 must come one cycle earlier than the others.
  
  "pathLatency": 6,
*/

/*
// Try to get a new output each clock cycle after an initially latency of 6. - ATTEMPT 1
// THIS DOESN'T WORK. Tries to put each input 'block' in a single data in stream. Due to different path latencies in the 2x2 conv tree,
//      input 'blocks' start mixing to give wrong output.
dataIn = {
16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
K2[15:0],L2in[175:160],16'd0,   K2[47:32],L2in[239:224],16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
K2[31:16],L2in[191:176],16'd0,  K2[63:48],L2in[255:240],16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0};
#2

dataIn = {
16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
K2[15:0],L2in[143:128],16'd0,   K2[47:32],L2in[207:192],16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
K2[31:16],L2in[159:144],16'd0,  K2[63:48],L2in[223:208],16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0};
#2

dataIn = {
16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
K2[15:0],L2in[47:32],16'd0,     K2[47:32],L2in[111:96],16'd0,   16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
K2[31:16],L2in[63:48],16'd0,    K2[63:48],L2in[127:112],16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0};
#2

dataIn = {
16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
K2[15:0],L2in[15:0],16'd0,     K2[47:32],L2in[79:64],16'd0,   16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
K2[31:16],L2in[31:16],16'd0,    K2[63:48],L2in[95:80],16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0};
#4
*/


// Try to get a new output each clock cycle after an initially latency of 6. - ATTEMPT 2
// THIS ONE WORKS. LATENCY MEANS NEEDS TO COME LATER. E.G. IF IN1 HAS LATENCY 2 AND IN3 HAS LATENCY 1, IN1 SHOULD COME 1 CYCLE AFTER IN3.
/*
layer2 in: 
IN2 X
IN4 r1c2 (in1)
IN6 X
IN8 r2c2 (in1)
*/
dataIn = {
16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
K2[15:0],L2in[175:160],16'd0,   K2[47:32],L2in[239:224],16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
K2[31:16],16'd0,16'd0,          K2[63:48],16'd0,16'd0,          16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0};
#2

/*
layer2 in: 
IN2 r1c1(in1)
IN4 r1c4 (in2)
IN6 r2c1(in1)
IN8 r2c4 (in2)
*/
dataIn = {
16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
K2[15:0],L2in[143:128],16'd0,   K2[47:32],L2in[207:192],16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
K2[31:16],L2in[191:176],16'd0,  K2[63:48],L2in[255:240],16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0};
#2

/*
layer2 in: 
IN2 r1c3(in2)
IN4 r3c2 (in3)
IN6 r2c3(in2)
IN8 r4c2 (in3)
*/
dataIn = {
16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
K2[15:0],L2in[47:32],16'd0,     K2[47:32],L2in[111:96],16'd0,   16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
K2[31:16],L2in[159:144],16'd0,  K2[63:48],L2in[223:208],16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0};
#2

/*
layer2 in: 
IN2 r3c1 (in3)
IN4 r3c4 (in4)
IN6 r4c1 (in3)
IN8 r4c4 (in4)
*/
dataIn = {
16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
K2[15:0],L2in[15:0],16'd0,      K2[47:32],L2in[79:64],16'd0,    16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
K2[31:16],L2in[63:48],16'd0,    K2[63:48],L2in[127:112],16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0};
#2

/*
layer2 in: 
IN2 r3c3 (in4)
IN4 X
IN6 r4c3 (in4)
IN8 X
*/
dataIn = {
16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
K2[15:0],16'd0,16'd0,           K2[47:32],16'd0,16'd0,          16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
K2[31:16],L2in[31:16],16'd0,    K2[63:48],L2in[95:80],16'd0,    16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  
16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,              16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0,  16'd0,16'd0,16'd0};
#2

dataIn = {16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0,16'd0};



end


endmodule